class transaction; 
  rand bit [15:0] A; 
  rand bit Load; 
  rand bit Left; 
  rand bit Din; 
  bit [15:0] register; 
  bit Dout; 
endclass:transaction
